//***************************************************************************************
//Ethernet packet class package
//This package include all the data members of the packet class
//***************************************************************************************

package Ethernet_packet_package;

`include "Ethernet_packet.sv"

endpackage: Ethernet_packet_package
